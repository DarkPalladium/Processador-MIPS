//Nomes:
//Pablo Miranda Batista 3482
//Roniel Nunes Barbosa 3464
//Samuel Aparecido D. Rodrigues 3476

module memoria(clk, memwrite, memread, memtoreg, aluresult, valor2, valorsalvar);
  input wire memwrite, memread, memtoreg, clk;
  input wire [31:0] aluresult, valor2;
  output reg [31:0] valorsalvar;

  reg [31:0] memorias [39:0];   //banco de Memoria


  initial begin
      memorias[0] = 32'b00000000000000000000000000000100;//4
      memorias[1] = 32'b00000000000000000000000000001000;//8
      memorias[2] = 32'b00000000000000000000000000010000;//16
      memorias[3] = 32'b00000000000000000000000000100000;//32
      memorias[4] = 32'b00000000000000000000000001000000;//64
      memorias[5] = 32'b00000000000000000000000010000000;//128
      memorias[6] = 32'b00000000000000000000000100000000;//256
      memorias[7] = 32'b00000000000000000000001000000000;//512
      memorias[8] = 32'b00000000000000000000010000000000;//1024
      memorias[9] = 32'b00000000000000000000100000000000;//2048
      memorias[10] = 32'b00000000000000000010000000000000;//4096
      memorias[11] = 32'b00000000000000000100000000000000;//8192
      memorias[12] = 32'b00000000000000001000000000000000;//16384
      memorias[13] = 32'b00000000000000000000000000000010;//2
      memorias[14] = 32'b00000000000000010000000000000000;//32768
      memorias[15] = 32'b00000000000000100000000000000000;//65536
      memorias[16] = 32'b00000000000000000000000000010101;//21
      memorias[17] = 32'b00000000000000000000000100010000;//272
      memorias[18] = 32'b00000000000000000000000001000100;//68
      memorias[19] = 32'b00000000000000000000000000000001;//1
      memorias[20] = 32'b00000000000000000000000000001111;//15
      memorias[21] = 32'b00000000000000000000000001000001;//65
      memorias[22] = 32'b00000000000000000000000001010101;//85
      memorias[23] = 32'b00000000000000000000000000001100;//12
      memorias[24] = 32'b00000000000000000000000000000011;//3
      memorias[25] = 32'b00000000000000000000000000000101;//5
      memorias[26] = 32'b00000000000000000000000000000110;//6
      memorias[27] = 32'b00000000000000000000000000000111;//7
      memorias[28] = 32'b00000000000000000000000000001001;//9
      memorias[29] = 32'b00000000000000000000000000001010;//10
      memorias[30] = 32'b00000000000000000000000000001011;//11
      memorias[31] = 32'b00000000000000000000000000001101;//13
      memorias[32] = 32'b00000000000000000000000000001110;//14
      memorias[33] = 32'b00000000000000000000000000010001;//17
      memorias[34] = 32'b00000000000000000000000000010100;//20
      memorias[35] = 32'b00000000000000000000000000011001;//25
      memorias[36] = 32'b00000000000000000000000000011110;//30
      memorias[37] = 32'b00000000000000000000000000100100;//36
      memorias[38] = 32'b00000000000000000000000000100010;//34
      memorias[39] = 32'b00000000000000000000000001000100;//68
  end

  always @ ( posedge clk ) begin
    if (memwrite) begin
      memorias[aluresult] = valor2;
    end
    if (memtoreg & memread) begin
      valorsalvar = memorias[aluresult];
    end
    if (~memtoreg) begin
      valorsalvar = aluresult;
    end
  end
endmodule //memoriamemwrite, memread, aluresult, data2, readdata);
